// NOT gate (74LS04/05)
module v7404 (input pin1, pin3, pin5, pin9, pin11, pin13,
				  output pin2, pin4, pin6, pin8, pin10, pin12);

	assign pin2 = !(pin1);
	assign pin4 = !(pin3);
	assign pin6 = !(pin5);
	
	assign pin8 = !(pin9);
	assign pin10 = !(pin11);
	assign pin12 = !(pin13);
	
endmodule